interface intf(input logic clk,rst);
  logic i0;
  logic i1;
  logic sel;
  logic y;
endinterface